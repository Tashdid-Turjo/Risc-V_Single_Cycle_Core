module alu;

endmodule