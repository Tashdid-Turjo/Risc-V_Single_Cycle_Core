// this module connected with '5.0.main_decoder' file //

