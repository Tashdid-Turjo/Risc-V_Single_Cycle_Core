// Step3

module Sign_Extend (In, ImmExt);
    
    input [31:0] In; // There's nothing written in the pic, so gave a name In.
    output [31:0] ImmExt;

    // It means -> In[31] is by default == 1'b1. Then MSB's 31:12 bits will be either 1 or 0 & LSB's 11:0 will be In's 31:20's value.
    assign ImmExt = {In[31]} ? {{20{1'b1}}, {In[31:20]}} :
                               {{20{1'b0}}, {In[31:20]}};

endmodule